parent(alice, bob).
parent(alice, bill).
parent(bob, carol).
parent(carol, dennis).
parent(carol, david).

ancestor(X, Y) :- parent(X, Y).
ancestor(X, Y) :- ancestor(X, Z), ancestor(Z, Y).
family(X, Y) :- ancestor(X, Y).
family(X, Y) :- family(Y, X).

age(alice, 30.00).
age(alice, Age)?
age(bob, 40.500).
age(bob, Age)?
weight(bob, 100.567000).
weight(bob, Weight)?

details(X, Age, Address, Weight) :- age(X, Age), address(X, Address), weight(X, Weight).
details(bob, Age, Address, Weight)?


family(X, Y)?
family(alice, Y)?
family(alex, Y)?
ancestor(bob, Y)?
address(bob, "10 someplace, somewhere").
address(bob, Address)?
address(carol, '123 "somestreet", sometown').
address(carol, Address)?