parent(alice, bob).
parent(alice, bill).
parent(bob, carol).
parent(carol, dennis).
parent(carol, david).
age(alice, 3000).
age(bob, 40500).
weight(bob, 100567000).

ancestor(X, Y) :- parent(X, Y).
ancestor(X, Y) :- ancestor(X, Z), ancestor(Z, Y).
family(X, Y) :- ancestor(X, Y).
family(X, Y) :- family(Y, X).

details(X, Age, Address, Weight) :- age(X, Age), address(X, Address), weight(X, Weight).
details(bob, Age, Address, Weight)?


age(alice, Age)?
age(bob, Age)?
weight(bob, Weight)?
family(X, Y)?
family(alice, Y)?
family(alex, Y)?
ancestor(bob, Y)?

address(bob, Address)?
address(carol, Address)?