p(0).
q(0).

p(1) :- p(0), q(1).
q(1) :- p(0), q(0).
p(2) :- p(1), q(2).
q(2) :- p(1), q(1).
p(3) :- p(2), q(3).
q(3) :- p(2), q(2).
p(4) :- p(3), q(4).
q(4) :- p(3), q(3).
p(5) :- p(4), q(5).
q(5) :- p(4), q(4).
p(6) :- p(5), q(6).
q(6) :- p(5), q(5).
p(7) :- p(6), q(7).
q(7) :- p(6), q(6).
p(8) :- p(7), q(8).
q(8) :- p(7), q(7).
p(9) :- p(8), q(9).
q(9) :- p(8), q(8).
p(10) :- p(9), q(10).
q(10) :- p(9), q(9).