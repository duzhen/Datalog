edge(a, b),
edge(a, c).
edge(b, d).
edge(c, d), edge(c, d).
edge(d, e).
not edge(f, e).

path(X, Y) :- edge(X, Y),
path(X, Y) := path(X, Z), path(Z, Y).
#path(X, X) = not edge(X, X).

path(a, b)?
path(f, X), f == e ?
path(a, X), path(X, d)?
#edge(f, e).