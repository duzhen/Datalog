p(0).
p(1).
k(0).

%positive cycle
k(1) :- p(2).
p(2) :- q(2).
q(2) :- k(0).

p(1) :- k(2).
q(2) :- p(2).
k(2) :- q(0).

%negation with positive cycle
m(1) :- not n(0).
n(0) :- not k(1).

q(X)?
k(X)?
n(X)?
m(X)?