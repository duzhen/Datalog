p(0).
q(Y).

p(1) :- not p(0).
p(1) :- p(0), X == 0.
p(X) :- p(0), p(Y), p(X, Y, Z), p(1, 2, 3).
p_(X) :- p(0), p(Y), p(Y, Z), p(1, 2, 3).

not q(X)?