p(0).

%positive cycle
k(1) :- p(2).
p(2) :- q(2).
q(2) :- k(0).

m(1) :- not n(0).
n(0) :- not k(1).
% p->q->k

q(X)?
k(X)?