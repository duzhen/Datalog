p(0).
q(0).

p(1) :- p(0), q(1).
q(1) :- p(0), q(0).
p(2) :- p(1), q(2).
q(2) :- p(1), q(1).
p(3) :- p(2), q(3).
q(3) :- p(2), q(2).
p(4) :- p(3), q(4).
q(4) :- p(3), q(3).
p(5) :- p(4), q(5).
q(5) :- p(4), q(4).
p(6) :- p(5), q(6).
q(6) :- p(5), q(5).
p(7) :- p(6), q(7).
q(7) :- p(6), q(6).
p(8) :- p(7), q(8).
q(8) :- p(7), q(7).
p(9) :- p(8), q(9).
q(9) :- p(8), q(8).
p(10) :- p(9), q(10).
q(10) :- p(9), q(9).
p(11) :- p(10), q(11).
q(11) :- p(10), q(10).
p(12) :- p(11), q(12).
q(12) :- p(11), q(11).
p(13) :- p(12), q(13).
q(13) :- p(12), q(12).
p(14) :- p(13), q(14).
q(14) :- p(13), q(13).
p(15) :- p(14), q(15).
q(15) :- p(14), q(14).
p(16) :- p(15), q(16).
q(16) :- p(15), q(15).
p(17) :- p(16), q(17).
q(17) :- p(16), q(16).
p(18) :- p(17), q(18).
q(18) :- p(17), q(17).
p(19) :- p(18), q(19).
q(19) :- p(18), q(18).
p(20) :- p(19), q(20).
q(20) :- p(19), q(19).
p(21) :- p(20), q(21).
q(21) :- p(20), q(20).
p(22) :- p(21), q(22).
q(22) :- p(21), q(21).
p(23) :- p(22), q(23).
q(23) :- p(22), q(22).
p(24) :- p(23), q(24).
q(24) :- p(23), q(23).
p(25) :- p(24), q(25).
q(25) :- p(24), q(24).
p(26) :- p(25), q(26).
q(26) :- p(25), q(25).
p(27) :- p(26), q(27).
q(27) :- p(26), q(26).
p(28) :- p(27), q(28).
q(28) :- p(27), q(27).
p(29) :- p(28), q(29).
q(29) :- p(28), q(28).
p(30) :- p(29), q(30).
q(30) :- p(29), q(29).
p(31) :- p(30), q(31).
q(31) :- p(30), q(30).
p(32) :- p(31), q(32).
q(32) :- p(31), q(31).
p(33) :- p(32), q(33).
q(33) :- p(32), q(32).
p(34) :- p(33), q(34).
q(34) :- p(33), q(33).
p(35) :- p(34), q(35).
q(35) :- p(34), q(34).
p(36) :- p(35), q(36).
q(36) :- p(35), q(35).
p(37) :- p(36), q(37).
q(37) :- p(36), q(36).
p(38) :- p(37), q(38).
q(38) :- p(37), q(37).
p(39) :- p(38), q(39).
q(39) :- p(38), q(38).
p(40) :- p(39), q(40).
q(40) :- p(39), q(39).
p(41) :- p(40), q(41).
q(41) :- p(40), q(40).
p(42) :- p(41), q(42).
q(42) :- p(41), q(41).
p(43) :- p(42), q(43).
q(43) :- p(42), q(42).
p(44) :- p(43), q(44).
q(44) :- p(43), q(43).
p(45) :- p(44), q(45).
q(45) :- p(44), q(44).
p(46) :- p(45), q(46).
q(46) :- p(45), q(45).
p(47) :- p(46), q(47).
q(47) :- p(46), q(46).
p(48) :- p(47), q(48).
q(48) :- p(47), q(47).
p(49) :- p(48), q(49).
q(49) :- p(48), q(48).
p(50) :- p(49), q(50).
q(50) :- p(49), q(49).
p(51) :- p(50), q(51).
q(51) :- p(50), q(50).
p(52) :- p(51), q(52).
q(52) :- p(51), q(51).
p(53) :- p(52), q(53).
q(53) :- p(52), q(52).
p(54) :- p(53), q(54).
q(54) :- p(53), q(53).
p(55) :- p(54), q(55).
q(55) :- p(54), q(54).
p(56) :- p(55), q(56).
q(56) :- p(55), q(55).
p(57) :- p(56), q(57).
q(57) :- p(56), q(56).
p(58) :- p(57), q(58).
q(58) :- p(57), q(57).
p(59) :- p(58), q(59).
q(59) :- p(58), q(58).
p(60) :- p(59), q(60).
q(60) :- p(59), q(59).
p(61) :- p(60), q(61).
q(61) :- p(60), q(60).
p(62) :- p(61), q(62).
q(62) :- p(61), q(61).
p(63) :- p(62), q(63).
q(63) :- p(62), q(62).
p(64) :- p(63), q(64).
q(64) :- p(63), q(63).
p(65) :- p(64), q(65).
q(65) :- p(64), q(64).
p(66) :- p(65), q(66).
q(66) :- p(65), q(65).
p(67) :- p(66), q(67).
q(67) :- p(66), q(66).
p(68) :- p(67), q(68).
q(68) :- p(67), q(67).
p(69) :- p(68), q(69).
q(69) :- p(68), q(68).
p(70) :- p(69), q(70).
q(70) :- p(69), q(69).
p(71) :- p(70), q(71).
q(71) :- p(70), q(70).
p(72) :- p(71), q(72).
q(72) :- p(71), q(71).
p(73) :- p(72), q(73).
q(73) :- p(72), q(72).
p(74) :- p(73), q(74).
q(74) :- p(73), q(73).
p(75) :- p(74), q(75).
q(75) :- p(74), q(74).
p(76) :- p(75), q(76).
q(76) :- p(75), q(75).
p(77) :- p(76), q(77).
q(77) :- p(76), q(76).
p(78) :- p(77), q(78).
q(78) :- p(77), q(77).
p(79) :- p(78), q(79).
q(79) :- p(78), q(78).
p(80) :- p(79), q(80).
q(80) :- p(79), q(79).
p(81) :- p(80), q(81).
q(81) :- p(80), q(80).
p(82) :- p(81), q(82).
q(82) :- p(81), q(81).
p(83) :- p(82), q(83).
q(83) :- p(82), q(82).
p(84) :- p(83), q(84).
q(84) :- p(83), q(83).
p(85) :- p(84), q(85).
q(85) :- p(84), q(84).
p(86) :- p(85), q(86).
q(86) :- p(85), q(85).
p(87) :- p(86), q(87).
q(87) :- p(86), q(86).
p(88) :- p(87), q(88).
q(88) :- p(87), q(87).
p(89) :- p(88), q(89).
q(89) :- p(88), q(88).
p(90) :- p(89), q(90).
q(90) :- p(89), q(89).
p(91) :- p(90), q(91).
q(91) :- p(90), q(90).
p(92) :- p(91), q(92).
q(92) :- p(91), q(91).
p(93) :- p(92), q(93).
q(93) :- p(92), q(92).
p(94) :- p(93), q(94).
q(94) :- p(93), q(93).
p(95) :- p(94), q(95).
q(95) :- p(94), q(94).
p(96) :- p(95), q(96).
q(96) :- p(95), q(95).
p(97) :- p(96), q(97).
q(97) :- p(96), q(96).
p(98) :- p(97), q(98).
q(98) :- p(97), q(97).
p(99) :- p(98), q(99).
q(99) :- p(98), q(98).
p(100) :- p(99), q(100).
q(100) :- p(99), q(99).
p(101) :- p(100), q(101).
q(101) :- p(100), q(100).
p(102) :- p(101), q(102).
q(102) :- p(101), q(101).
p(103) :- p(102), q(103).
q(103) :- p(102), q(102).
p(104) :- p(103), q(104).
q(104) :- p(103), q(103).
p(105) :- p(104), q(105).
q(105) :- p(104), q(104).
p(106) :- p(105), q(106).
q(106) :- p(105), q(105).
p(107) :- p(106), q(107).
q(107) :- p(106), q(106).
p(108) :- p(107), q(108).
q(108) :- p(107), q(107).
p(109) :- p(108), q(109).
q(109) :- p(108), q(108).
p(110) :- p(109), q(110).
q(110) :- p(109), q(109).
p(111) :- p(110), q(111).
q(111) :- p(110), q(110).
p(112) :- p(111), q(112).
q(112) :- p(111), q(111).
p(113) :- p(112), q(113).
q(113) :- p(112), q(112).
p(114) :- p(113), q(114).
q(114) :- p(113), q(113).
p(115) :- p(114), q(115).
q(115) :- p(114), q(114).
p(116) :- p(115), q(116).
q(116) :- p(115), q(115).
p(117) :- p(116), q(117).
q(117) :- p(116), q(116).
p(118) :- p(117), q(118).
q(118) :- p(117), q(117).
p(119) :- p(118), q(119).
q(119) :- p(118), q(118).
p(120) :- p(119), q(120).
q(120) :- p(119), q(119).
p(121) :- p(120), q(121).
q(121) :- p(120), q(120).
p(122) :- p(121), q(122).
q(122) :- p(121), q(121).
p(123) :- p(122), q(123).
q(123) :- p(122), q(122).
p(124) :- p(123), q(124).
q(124) :- p(123), q(123).
p(125) :- p(124), q(125).
q(125) :- p(124), q(124).
p(126) :- p(125), q(126).
q(126) :- p(125), q(125).
p(127) :- p(126), q(127).
q(127) :- p(126), q(126).
p(128) :- p(127), q(128).
q(128) :- p(127), q(127).
p(129) :- p(128), q(129).
q(129) :- p(128), q(128).
p(130) :- p(129), q(130).
q(130) :- p(129), q(129).
p(131) :- p(130), q(131).
q(131) :- p(130), q(130).
p(132) :- p(131), q(132).
q(132) :- p(131), q(131).
p(133) :- p(132), q(133).
q(133) :- p(132), q(132).
p(134) :- p(133), q(134).
q(134) :- p(133), q(133).
p(135) :- p(134), q(135).
q(135) :- p(134), q(134).
p(136) :- p(135), q(136).
q(136) :- p(135), q(135).
p(137) :- p(136), q(137).
q(137) :- p(136), q(136).
p(138) :- p(137), q(138).
q(138) :- p(137), q(137).
p(139) :- p(138), q(139).
q(139) :- p(138), q(138).
p(140) :- p(139), q(140).
q(140) :- p(139), q(139).
p(141) :- p(140), q(141).
q(141) :- p(140), q(140).
p(142) :- p(141), q(142).
q(142) :- p(141), q(141).
p(143) :- p(142), q(143).
q(143) :- p(142), q(142).
p(144) :- p(143), q(144).
q(144) :- p(143), q(143).
p(145) :- p(144), q(145).
q(145) :- p(144), q(144).
p(146) :- p(145), q(146).
q(146) :- p(145), q(145).
p(147) :- p(146), q(147).
q(147) :- p(146), q(146).
p(148) :- p(147), q(148).
q(148) :- p(147), q(147).
p(149) :- p(148), q(149).
q(149) :- p(148), q(148).
p(150) :- p(149), q(150).
q(150) :- p(149), q(149).
p(151) :- p(150), q(151).
q(151) :- p(150), q(150).
p(152) :- p(151), q(152).
q(152) :- p(151), q(151).
p(153) :- p(152), q(153).
q(153) :- p(152), q(152).
p(154) :- p(153), q(154).
q(154) :- p(153), q(153).
p(155) :- p(154), q(155).
q(155) :- p(154), q(154).
p(156) :- p(155), q(156).
q(156) :- p(155), q(155).
p(157) :- p(156), q(157).
q(157) :- p(156), q(156).
p(158) :- p(157), q(158).
q(158) :- p(157), q(157).
p(159) :- p(158), q(159).
q(159) :- p(158), q(158).
p(160) :- p(159), q(160).
q(160) :- p(159), q(159).
p(161) :- p(160), q(161).
q(161) :- p(160), q(160).
p(162) :- p(161), q(162).
q(162) :- p(161), q(161).
p(163) :- p(162), q(163).
q(163) :- p(162), q(162).
p(164) :- p(163), q(164).
q(164) :- p(163), q(163).
p(165) :- p(164), q(165).
q(165) :- p(164), q(164).
p(166) :- p(165), q(166).
q(166) :- p(165), q(165).
p(167) :- p(166), q(167).
q(167) :- p(166), q(166).
p(168) :- p(167), q(168).
q(168) :- p(167), q(167).
p(169) :- p(168), q(169).
q(169) :- p(168), q(168).
p(170) :- p(169), q(170).
q(170) :- p(169), q(169).
p(171) :- p(170), q(171).
q(171) :- p(170), q(170).
p(172) :- p(171), q(172).
q(172) :- p(171), q(171).
p(173) :- p(172), q(173).
q(173) :- p(172), q(172).
p(174) :- p(173), q(174).
q(174) :- p(173), q(173).
p(175) :- p(174), q(175).
q(175) :- p(174), q(174).
p(176) :- p(175), q(176).
q(176) :- p(175), q(175).
p(177) :- p(176), q(177).
q(177) :- p(176), q(176).
p(178) :- p(177), q(178).
q(178) :- p(177), q(177).
p(179) :- p(178), q(179).
q(179) :- p(178), q(178).
p(180) :- p(179), q(180).
q(180) :- p(179), q(179).
p(181) :- p(180), q(181).
q(181) :- p(180), q(180).
p(182) :- p(181), q(182).
q(182) :- p(181), q(181).
p(183) :- p(182), q(183).
q(183) :- p(182), q(182).
p(184) :- p(183), q(184).
q(184) :- p(183), q(183).
p(185) :- p(184), q(185).
q(185) :- p(184), q(184).
p(186) :- p(185), q(186).
q(186) :- p(185), q(185).
p(187) :- p(186), q(187).
q(187) :- p(186), q(186).
p(188) :- p(187), q(188).
q(188) :- p(187), q(187).
p(189) :- p(188), q(189).
q(189) :- p(188), q(188).
p(190) :- p(189), q(190).
q(190) :- p(189), q(189).
p(191) :- p(190), q(191).
q(191) :- p(190), q(190).
p(192) :- p(191), q(192).
q(192) :- p(191), q(191).
p(193) :- p(192), q(193).
q(193) :- p(192), q(192).
p(194) :- p(193), q(194).
q(194) :- p(193), q(193).
p(195) :- p(194), q(195).
q(195) :- p(194), q(194).
p(196) :- p(195), q(196).
q(196) :- p(195), q(195).
p(197) :- p(196), q(197).
q(197) :- p(196), q(196).
p(198) :- p(197), q(198).
q(198) :- p(197), q(197).
p(199) :- p(198), q(199).
q(199) :- p(198), q(198).
p(200) :- p(199), q(200).
q(200) :- p(199), q(199).
p(201) :- p(200), q(201).
q(201) :- p(200), q(200).
p(202) :- p(201), q(202).
q(202) :- p(201), q(201).
p(203) :- p(202), q(203).
q(203) :- p(202), q(202).
p(204) :- p(203), q(204).
q(204) :- p(203), q(203).
p(205) :- p(204), q(205).
q(205) :- p(204), q(204).
p(206) :- p(205), q(206).
q(206) :- p(205), q(205).
p(207) :- p(206), q(207).
q(207) :- p(206), q(206).
p(208) :- p(207), q(208).
q(208) :- p(207), q(207).
p(209) :- p(208), q(209).
q(209) :- p(208), q(208).
p(210) :- p(209), q(210).
q(210) :- p(209), q(209).
p(211) :- p(210), q(211).
q(211) :- p(210), q(210).
p(212) :- p(211), q(212).
q(212) :- p(211), q(211).
p(213) :- p(212), q(213).
q(213) :- p(212), q(212).
p(214) :- p(213), q(214).
q(214) :- p(213), q(213).
p(215) :- p(214), q(215).
q(215) :- p(214), q(214).
p(216) :- p(215), q(216).
q(216) :- p(215), q(215).
p(217) :- p(216), q(217).
q(217) :- p(216), q(216).
p(218) :- p(217), q(218).
q(218) :- p(217), q(217).
p(219) :- p(218), q(219).
q(219) :- p(218), q(218).
p(220) :- p(219), q(220).
q(220) :- p(219), q(219).
p(221) :- p(220), q(221).
q(221) :- p(220), q(220).
p(222) :- p(221), q(222).
q(222) :- p(221), q(221).
p(223) :- p(222), q(223).
q(223) :- p(222), q(222).
p(224) :- p(223), q(224).
q(224) :- p(223), q(223).
p(225) :- p(224), q(225).
q(225) :- p(224), q(224).
p(226) :- p(225), q(226).
q(226) :- p(225), q(225).
p(227) :- p(226), q(227).
q(227) :- p(226), q(226).
p(228) :- p(227), q(228).
q(228) :- p(227), q(227).
p(229) :- p(228), q(229).
q(229) :- p(228), q(228).
p(230) :- p(229), q(230).
q(230) :- p(229), q(229).
p(231) :- p(230), q(231).
q(231) :- p(230), q(230).
p(232) :- p(231), q(232).
q(232) :- p(231), q(231).
p(233) :- p(232), q(233).
q(233) :- p(232), q(232).
p(234) :- p(233), q(234).
q(234) :- p(233), q(233).
p(235) :- p(234), q(235).
q(235) :- p(234), q(234).
p(236) :- p(235), q(236).
q(236) :- p(235), q(235).
p(237) :- p(236), q(237).
q(237) :- p(236), q(236).
p(238) :- p(237), q(238).
q(238) :- p(237), q(237).
p(239) :- p(238), q(239).
q(239) :- p(238), q(238).
p(240) :- p(239), q(240).
q(240) :- p(239), q(239).
p(241) :- p(240), q(241).
q(241) :- p(240), q(240).
p(242) :- p(241), q(242).
q(242) :- p(241), q(241).
p(243) :- p(242), q(243).
q(243) :- p(242), q(242).
p(244) :- p(243), q(244).
q(244) :- p(243), q(243).
p(245) :- p(244), q(245).
q(245) :- p(244), q(244).
p(246) :- p(245), q(246).
q(246) :- p(245), q(245).
p(247) :- p(246), q(247).
q(247) :- p(246), q(246).
p(248) :- p(247), q(248).
q(248) :- p(247), q(247).
p(249) :- p(248), q(249).
q(249) :- p(248), q(248).
p(250) :- p(249), q(250).
q(250) :- p(249), q(249).
p(251) :- p(250), q(251).
q(251) :- p(250), q(250).
p(252) :- p(251), q(252).
q(252) :- p(251), q(251).
p(253) :- p(252), q(253).
q(253) :- p(252), q(252).
p(254) :- p(253), q(254).
q(254) :- p(253), q(253).
p(255) :- p(254), q(255).
q(255) :- p(254), q(254).
p(256) :- p(255), q(256).
q(256) :- p(255), q(255).
p(257) :- p(256), q(257).
q(257) :- p(256), q(256).
p(258) :- p(257), q(258).
q(258) :- p(257), q(257).
p(259) :- p(258), q(259).
q(259) :- p(258), q(258).
p(260) :- p(259), q(260).
q(260) :- p(259), q(259).
p(261) :- p(260), q(261).
q(261) :- p(260), q(260).
p(262) :- p(261), q(262).
q(262) :- p(261), q(261).
p(263) :- p(262), q(263).
q(263) :- p(262), q(262).
p(264) :- p(263), q(264).
q(264) :- p(263), q(263).
p(265) :- p(264), q(265).
q(265) :- p(264), q(264).
p(266) :- p(265), q(266).
q(266) :- p(265), q(265).
p(267) :- p(266), q(267).
q(267) :- p(266), q(266).
p(268) :- p(267), q(268).
q(268) :- p(267), q(267).
p(269) :- p(268), q(269).
q(269) :- p(268), q(268).
p(270) :- p(269), q(270).
q(270) :- p(269), q(269).
p(271) :- p(270), q(271).
q(271) :- p(270), q(270).
p(272) :- p(271), q(272).
q(272) :- p(271), q(271).
p(273) :- p(272), q(273).
q(273) :- p(272), q(272).
p(274) :- p(273), q(274).
q(274) :- p(273), q(273).
p(275) :- p(274), q(275).
q(275) :- p(274), q(274).
p(276) :- p(275), q(276).
q(276) :- p(275), q(275).
p(277) :- p(276), q(277).
q(277) :- p(276), q(276).
p(278) :- p(277), q(278).
q(278) :- p(277), q(277).
p(279) :- p(278), q(279).
q(279) :- p(278), q(278).
p(280) :- p(279), q(280).
q(280) :- p(279), q(279).
p(281) :- p(280), q(281).
q(281) :- p(280), q(280).
p(282) :- p(281), q(282).
q(282) :- p(281), q(281).
p(283) :- p(282), q(283).
q(283) :- p(282), q(282).
p(284) :- p(283), q(284).
q(284) :- p(283), q(283).
p(285) :- p(284), q(285).
q(285) :- p(284), q(284).
p(286) :- p(285), q(286).
q(286) :- p(285), q(285).
p(287) :- p(286), q(287).
q(287) :- p(286), q(286).
p(288) :- p(287), q(288).
q(288) :- p(287), q(287).
p(289) :- p(288), q(289).
q(289) :- p(288), q(288).
p(290) :- p(289), q(290).
q(290) :- p(289), q(289).
p(291) :- p(290), q(291).
q(291) :- p(290), q(290).
p(292) :- p(291), q(292).
q(292) :- p(291), q(291).
p(293) :- p(292), q(293).
q(293) :- p(292), q(292).
p(294) :- p(293), q(294).
q(294) :- p(293), q(293).
p(295) :- p(294), q(295).
q(295) :- p(294), q(294).
p(296) :- p(295), q(296).
q(296) :- p(295), q(295).
p(297) :- p(296), q(297).
q(297) :- p(296), q(296).
p(298) :- p(297), q(298).
q(298) :- p(297), q(297).
p(299) :- p(298), q(299).
q(299) :- p(298), q(298).
p(300) :- p(299), q(300).
q(300) :- p(299), q(299).
p(301) :- p(300), q(301).
q(301) :- p(300), q(300).
p(302) :- p(301), q(302).
q(302) :- p(301), q(301).
p(303) :- p(302), q(303).
q(303) :- p(302), q(302).
p(304) :- p(303), q(304).
q(304) :- p(303), q(303).
p(305) :- p(304), q(305).
q(305) :- p(304), q(304).
p(306) :- p(305), q(306).
q(306) :- p(305), q(305).
p(307) :- p(306), q(307).
q(307) :- p(306), q(306).
p(308) :- p(307), q(308).
q(308) :- p(307), q(307).
p(309) :- p(308), q(309).
q(309) :- p(308), q(308).
p(310) :- p(309), q(310).
q(310) :- p(309), q(309).
p(311) :- p(310), q(311).
q(311) :- p(310), q(310).
p(312) :- p(311), q(312).
q(312) :- p(311), q(311).
p(313) :- p(312), q(313).
q(313) :- p(312), q(312).
p(314) :- p(313), q(314).
q(314) :- p(313), q(313).
p(315) :- p(314), q(315).
q(315) :- p(314), q(314).
p(316) :- p(315), q(316).
q(316) :- p(315), q(315).
p(317) :- p(316), q(317).
q(317) :- p(316), q(316).
p(318) :- p(317), q(318).
q(318) :- p(317), q(317).
p(319) :- p(318), q(319).
q(319) :- p(318), q(318).
p(320) :- p(319), q(320).
q(320) :- p(319), q(319).
p(321) :- p(320), q(321).
q(321) :- p(320), q(320).
p(322) :- p(321), q(322).
q(322) :- p(321), q(321).
p(323) :- p(322), q(323).
q(323) :- p(322), q(322).
p(324) :- p(323), q(324).
q(324) :- p(323), q(323).
p(325) :- p(324), q(325).
q(325) :- p(324), q(324).
p(326) :- p(325), q(326).
q(326) :- p(325), q(325).
p(327) :- p(326), q(327).
q(327) :- p(326), q(326).
p(328) :- p(327), q(328).
q(328) :- p(327), q(327).
p(329) :- p(328), q(329).
q(329) :- p(328), q(328).
p(330) :- p(329), q(330).
q(330) :- p(329), q(329).
p(331) :- p(330), q(331).
q(331) :- p(330), q(330).
p(332) :- p(331), q(332).
q(332) :- p(331), q(331).
p(333) :- p(332), q(333).
q(333) :- p(332), q(332).
p(334) :- p(333), q(334).
q(334) :- p(333), q(333).
p(335) :- p(334), q(335).
q(335) :- p(334), q(334).
p(336) :- p(335), q(336).
q(336) :- p(335), q(335).
p(337) :- p(336), q(337).
q(337) :- p(336), q(336).
p(338) :- p(337), q(338).
q(338) :- p(337), q(337).
p(339) :- p(338), q(339).
q(339) :- p(338), q(338).
p(340) :- p(339), q(340).
q(340) :- p(339), q(339).
p(341) :- p(340), q(341).
q(341) :- p(340), q(340).
p(342) :- p(341), q(342).
q(342) :- p(341), q(341).
p(343) :- p(342), q(343).
q(343) :- p(342), q(342).
p(344) :- p(343), q(344).
q(344) :- p(343), q(343).
p(345) :- p(344), q(345).
q(345) :- p(344), q(344).
p(346) :- p(345), q(346).
q(346) :- p(345), q(345).
p(347) :- p(346), q(347).
q(347) :- p(346), q(346).
p(348) :- p(347), q(348).
q(348) :- p(347), q(347).
p(349) :- p(348), q(349).
q(349) :- p(348), q(348).
p(350) :- p(349), q(350).
q(350) :- p(349), q(349).
p(351) :- p(350), q(351).
q(351) :- p(350), q(350).
p(352) :- p(351), q(352).
q(352) :- p(351), q(351).
p(353) :- p(352), q(353).
q(353) :- p(352), q(352).
p(354) :- p(353), q(354).
q(354) :- p(353), q(353).
p(355) :- p(354), q(355).
q(355) :- p(354), q(354).
p(356) :- p(355), q(356).
q(356) :- p(355), q(355).
p(357) :- p(356), q(357).
q(357) :- p(356), q(356).
p(358) :- p(357), q(358).
q(358) :- p(357), q(357).
p(359) :- p(358), q(359).
q(359) :- p(358), q(358).
p(360) :- p(359), q(360).
q(360) :- p(359), q(359).
p(361) :- p(360), q(361).
q(361) :- p(360), q(360).
p(362) :- p(361), q(362).
q(362) :- p(361), q(361).
p(363) :- p(362), q(363).
q(363) :- p(362), q(362).
p(364) :- p(363), q(364).
q(364) :- p(363), q(363).
p(365) :- p(364), q(365).
q(365) :- p(364), q(364).
p(366) :- p(365), q(366).
q(366) :- p(365), q(365).
p(367) :- p(366), q(367).
q(367) :- p(366), q(366).
p(368) :- p(367), q(368).
q(368) :- p(367), q(367).
p(369) :- p(368), q(369).
q(369) :- p(368), q(368).
p(370) :- p(369), q(370).
q(370) :- p(369), q(369).
p(371) :- p(370), q(371).
q(371) :- p(370), q(370).
p(372) :- p(371), q(372).
q(372) :- p(371), q(371).
p(373) :- p(372), q(373).
q(373) :- p(372), q(372).
p(374) :- p(373), q(374).
q(374) :- p(373), q(373).
p(375) :- p(374), q(375).
q(375) :- p(374), q(374).
p(376) :- p(375), q(376).
q(376) :- p(375), q(375).
p(377) :- p(376), q(377).
q(377) :- p(376), q(376).
p(378) :- p(377), q(378).
q(378) :- p(377), q(377).
p(379) :- p(378), q(379).
q(379) :- p(378), q(378).
p(380) :- p(379), q(380).
q(380) :- p(379), q(379).
p(381) :- p(380), q(381).
q(381) :- p(380), q(380).
p(382) :- p(381), q(382).
q(382) :- p(381), q(381).
p(383) :- p(382), q(383).
q(383) :- p(382), q(382).
p(384) :- p(383), q(384).
q(384) :- p(383), q(383).
p(385) :- p(384), q(385).
q(385) :- p(384), q(384).
p(386) :- p(385), q(386).
q(386) :- p(385), q(385).
p(387) :- p(386), q(387).
q(387) :- p(386), q(386).
p(388) :- p(387), q(388).
q(388) :- p(387), q(387).
p(389) :- p(388), q(389).
q(389) :- p(388), q(388).
p(390) :- p(389), q(390).
q(390) :- p(389), q(389).
p(391) :- p(390), q(391).
q(391) :- p(390), q(390).
p(392) :- p(391), q(392).
q(392) :- p(391), q(391).
p(393) :- p(392), q(393).
q(393) :- p(392), q(392).
p(394) :- p(393), q(394).
q(394) :- p(393), q(393).
p(395) :- p(394), q(395).
q(395) :- p(394), q(394).
p(396) :- p(395), q(396).
q(396) :- p(395), q(395).
p(397) :- p(396), q(397).
q(397) :- p(396), q(396).
p(398) :- p(397), q(398).
q(398) :- p(397), q(397).
p(399) :- p(398), q(399).
q(399) :- p(398), q(398).
p(400) :- p(399), q(400).
q(400) :- p(399), q(399).
p(401) :- p(400), q(401).
q(401) :- p(400), q(400).
p(402) :- p(401), q(402).
q(402) :- p(401), q(401).
p(403) :- p(402), q(403).
q(403) :- p(402), q(402).
p(404) :- p(403), q(404).
q(404) :- p(403), q(403).
p(405) :- p(404), q(405).
q(405) :- p(404), q(404).
p(406) :- p(405), q(406).
q(406) :- p(405), q(405).
p(407) :- p(406), q(407).
q(407) :- p(406), q(406).
p(408) :- p(407), q(408).
q(408) :- p(407), q(407).
p(409) :- p(408), q(409).
q(409) :- p(408), q(408).
p(410) :- p(409), q(410).
q(410) :- p(409), q(409).
p(411) :- p(410), q(411).
q(411) :- p(410), q(410).
p(412) :- p(411), q(412).
q(412) :- p(411), q(411).
p(413) :- p(412), q(413).
q(413) :- p(412), q(412).
p(414) :- p(413), q(414).
q(414) :- p(413), q(413).
p(415) :- p(414), q(415).
q(415) :- p(414), q(414).
p(416) :- p(415), q(416).
q(416) :- p(415), q(415).
p(417) :- p(416), q(417).
q(417) :- p(416), q(416).
p(418) :- p(417), q(418).
q(418) :- p(417), q(417).
p(419) :- p(418), q(419).
q(419) :- p(418), q(418).
p(420) :- p(419), q(420).
q(420) :- p(419), q(419).
p(421) :- p(420), q(421).
q(421) :- p(420), q(420).
p(422) :- p(421), q(422).
q(422) :- p(421), q(421).
p(423) :- p(422), q(423).
q(423) :- p(422), q(422).
p(424) :- p(423), q(424).
q(424) :- p(423), q(423).
p(425) :- p(424), q(425).
q(425) :- p(424), q(424).
p(426) :- p(425), q(426).
q(426) :- p(425), q(425).
p(427) :- p(426), q(427).
q(427) :- p(426), q(426).
p(428) :- p(427), q(428).
q(428) :- p(427), q(427).
p(429) :- p(428), q(429).
q(429) :- p(428), q(428).
p(430) :- p(429), q(430).
q(430) :- p(429), q(429).
p(431) :- p(430), q(431).
q(431) :- p(430), q(430).
p(432) :- p(431), q(432).
q(432) :- p(431), q(431).
p(433) :- p(432), q(433).
q(433) :- p(432), q(432).
p(434) :- p(433), q(434).
q(434) :- p(433), q(433).
p(435) :- p(434), q(435).
q(435) :- p(434), q(434).
p(436) :- p(435), q(436).
q(436) :- p(435), q(435).
p(437) :- p(436), q(437).
q(437) :- p(436), q(436).
p(438) :- p(437), q(438).
q(438) :- p(437), q(437).
p(439) :- p(438), q(439).
q(439) :- p(438), q(438).
p(440) :- p(439), q(440).
q(440) :- p(439), q(439).
p(441) :- p(440), q(441).
q(441) :- p(440), q(440).
p(442) :- p(441), q(442).
q(442) :- p(441), q(441).
p(443) :- p(442), q(443).
q(443) :- p(442), q(442).
p(444) :- p(443), q(444).
q(444) :- p(443), q(443).
p(445) :- p(444), q(445).
q(445) :- p(444), q(444).
p(446) :- p(445), q(446).
q(446) :- p(445), q(445).
p(447) :- p(446), q(447).
q(447) :- p(446), q(446).
p(448) :- p(447), q(448).
q(448) :- p(447), q(447).
p(449) :- p(448), q(449).
q(449) :- p(448), q(448).
p(450) :- p(449), q(450).
q(450) :- p(449), q(449).
p(451) :- p(450), q(451).
q(451) :- p(450), q(450).
p(452) :- p(451), q(452).
q(452) :- p(451), q(451).
p(453) :- p(452), q(453).
q(453) :- p(452), q(452).
p(454) :- p(453), q(454).
q(454) :- p(453), q(453).
p(455) :- p(454), q(455).
q(455) :- p(454), q(454).
p(456) :- p(455), q(456).
q(456) :- p(455), q(455).
p(457) :- p(456), q(457).
q(457) :- p(456), q(456).
p(458) :- p(457), q(458).
q(458) :- p(457), q(457).
p(459) :- p(458), q(459).
q(459) :- p(458), q(458).
p(460) :- p(459), q(460).
q(460) :- p(459), q(459).
p(461) :- p(460), q(461).
q(461) :- p(460), q(460).
p(462) :- p(461), q(462).
q(462) :- p(461), q(461).
p(463) :- p(462), q(463).
q(463) :- p(462), q(462).
p(464) :- p(463), q(464).
q(464) :- p(463), q(463).
p(465) :- p(464), q(465).
q(465) :- p(464), q(464).
p(466) :- p(465), q(466).
q(466) :- p(465), q(465).
p(467) :- p(466), q(467).
q(467) :- p(466), q(466).
p(468) :- p(467), q(468).
q(468) :- p(467), q(467).
p(469) :- p(468), q(469).
q(469) :- p(468), q(468).
p(470) :- p(469), q(470).
q(470) :- p(469), q(469).
p(471) :- p(470), q(471).
q(471) :- p(470), q(470).
p(472) :- p(471), q(472).
q(472) :- p(471), q(471).
p(473) :- p(472), q(473).
q(473) :- p(472), q(472).
p(474) :- p(473), q(474).
q(474) :- p(473), q(473).
p(475) :- p(474), q(475).
q(475) :- p(474), q(474).
p(476) :- p(475), q(476).
q(476) :- p(475), q(475).
p(477) :- p(476), q(477).
q(477) :- p(476), q(476).
p(478) :- p(477), q(478).
q(478) :- p(477), q(477).
p(479) :- p(478), q(479).
q(479) :- p(478), q(478).
p(480) :- p(479), q(480).
q(480) :- p(479), q(479).
p(481) :- p(480), q(481).
q(481) :- p(480), q(480).
p(482) :- p(481), q(482).
q(482) :- p(481), q(481).
p(483) :- p(482), q(483).
q(483) :- p(482), q(482).
p(484) :- p(483), q(484).
q(484) :- p(483), q(483).
p(485) :- p(484), q(485).
q(485) :- p(484), q(484).
p(486) :- p(485), q(486).
q(486) :- p(485), q(485).
p(487) :- p(486), q(487).
q(487) :- p(486), q(486).
p(488) :- p(487), q(488).
q(488) :- p(487), q(487).
p(489) :- p(488), q(489).
q(489) :- p(488), q(488).
p(490) :- p(489), q(490).
q(490) :- p(489), q(489).
p(491) :- p(490), q(491).
q(491) :- p(490), q(490).
p(492) :- p(491), q(492).
q(492) :- p(491), q(491).
p(493) :- p(492), q(493).
q(493) :- p(492), q(492).
p(494) :- p(493), q(494).
q(494) :- p(493), q(493).
p(495) :- p(494), q(495).
q(495) :- p(494), q(494).
p(496) :- p(495), q(496).
q(496) :- p(495), q(495).
p(497) :- p(496), q(497).
q(497) :- p(496), q(496).
p(498) :- p(497), q(498).
q(498) :- p(497), q(497).
p(499) :- p(498), q(499).
q(499) :- p(498), q(498).
p(500) :- p(499), q(500).
q(500) :- p(499), q(499).
p(501) :- p(500), q(501).
q(501) :- p(500), q(500).
p(502) :- p(501), q(502).
q(502) :- p(501), q(501).
p(503) :- p(502), q(503).
q(503) :- p(502), q(502).
p(504) :- p(503), q(504).
q(504) :- p(503), q(503).
p(505) :- p(504), q(505).
q(505) :- p(504), q(504).
p(506) :- p(505), q(506).
q(506) :- p(505), q(505).
p(507) :- p(506), q(507).
q(507) :- p(506), q(506).
p(508) :- p(507), q(508).
q(508) :- p(507), q(507).
p(509) :- p(508), q(509).
q(509) :- p(508), q(508).
p(510) :- p(509), q(510).
q(510) :- p(509), q(509).
p(511) :- p(510), q(511).
q(511) :- p(510), q(510).
p(512) :- p(511), q(512).
q(512) :- p(511), q(511).
p(513) :- p(512), q(513).
q(513) :- p(512), q(512).
p(514) :- p(513), q(514).
q(514) :- p(513), q(513).
p(515) :- p(514), q(515).
q(515) :- p(514), q(514).
p(516) :- p(515), q(516).
q(516) :- p(515), q(515).
p(517) :- p(516), q(517).
q(517) :- p(516), q(516).
p(518) :- p(517), q(518).
q(518) :- p(517), q(517).
p(519) :- p(518), q(519).
q(519) :- p(518), q(518).
p(520) :- p(519), q(520).
q(520) :- p(519), q(519).
p(521) :- p(520), q(521).
q(521) :- p(520), q(520).
p(522) :- p(521), q(522).
q(522) :- p(521), q(521).
p(523) :- p(522), q(523).
q(523) :- p(522), q(522).
p(524) :- p(523), q(524).
q(524) :- p(523), q(523).
p(525) :- p(524), q(525).
q(525) :- p(524), q(524).
p(526) :- p(525), q(526).
q(526) :- p(525), q(525).
p(527) :- p(526), q(527).
q(527) :- p(526), q(526).
p(528) :- p(527), q(528).
q(528) :- p(527), q(527).
p(529) :- p(528), q(529).
q(529) :- p(528), q(528).
p(530) :- p(529), q(530).
q(530) :- p(529), q(529).
p(531) :- p(530), q(531).
q(531) :- p(530), q(530).
p(532) :- p(531), q(532).
q(532) :- p(531), q(531).
p(533) :- p(532), q(533).
q(533) :- p(532), q(532).
p(534) :- p(533), q(534).
q(534) :- p(533), q(533).
p(535) :- p(534), q(535).
q(535) :- p(534), q(534).
p(536) :- p(535), q(536).
q(536) :- p(535), q(535).
p(537) :- p(536), q(537).
q(537) :- p(536), q(536).
p(538) :- p(537), q(538).
q(538) :- p(537), q(537).
p(539) :- p(538), q(539).
q(539) :- p(538), q(538).
p(540) :- p(539), q(540).
q(540) :- p(539), q(539).
p(541) :- p(540), q(541).
q(541) :- p(540), q(540).
p(542) :- p(541), q(542).
q(542) :- p(541), q(541).
p(543) :- p(542), q(543).
q(543) :- p(542), q(542).
p(544) :- p(543), q(544).
q(544) :- p(543), q(543).
p(545) :- p(544), q(545).
q(545) :- p(544), q(544).
p(546) :- p(545), q(546).
q(546) :- p(545), q(545).
p(547) :- p(546), q(547).
q(547) :- p(546), q(546).
p(548) :- p(547), q(548).
q(548) :- p(547), q(547).
p(549) :- p(548), q(549).
q(549) :- p(548), q(548).
p(550) :- p(549), q(550).
q(550) :- p(549), q(549).
p(551) :- p(550), q(551).
q(551) :- p(550), q(550).
p(552) :- p(551), q(552).
q(552) :- p(551), q(551).
p(553) :- p(552), q(553).
q(553) :- p(552), q(552).
p(554) :- p(553), q(554).
q(554) :- p(553), q(553).
p(555) :- p(554), q(555).
q(555) :- p(554), q(554).
p(556) :- p(555), q(556).
q(556) :- p(555), q(555).
p(557) :- p(556), q(557).
q(557) :- p(556), q(556).
p(558) :- p(557), q(558).
q(558) :- p(557), q(557).
p(559) :- p(558), q(559).
q(559) :- p(558), q(558).
p(560) :- p(559), q(560).
q(560) :- p(559), q(559).
p(561) :- p(560), q(561).
q(561) :- p(560), q(560).
p(562) :- p(561), q(562).
q(562) :- p(561), q(561).
p(563) :- p(562), q(563).
q(563) :- p(562), q(562).
p(564) :- p(563), q(564).
q(564) :- p(563), q(563).
p(565) :- p(564), q(565).
q(565) :- p(564), q(564).
p(566) :- p(565), q(566).
q(566) :- p(565), q(565).
p(567) :- p(566), q(567).
q(567) :- p(566), q(566).
p(568) :- p(567), q(568).
q(568) :- p(567), q(567).
p(569) :- p(568), q(569).
q(569) :- p(568), q(568).
p(570) :- p(569), q(570).
q(570) :- p(569), q(569).
p(571) :- p(570), q(571).
q(571) :- p(570), q(570).
p(572) :- p(571), q(572).
q(572) :- p(571), q(571).
p(573) :- p(572), q(573).
q(573) :- p(572), q(572).
p(574) :- p(573), q(574).
q(574) :- p(573), q(573).
p(575) :- p(574), q(575).
q(575) :- p(574), q(574).
p(576) :- p(575), q(576).
q(576) :- p(575), q(575).
p(577) :- p(576), q(577).
q(577) :- p(576), q(576).
p(578) :- p(577), q(578).
q(578) :- p(577), q(577).
p(579) :- p(578), q(579).
q(579) :- p(578), q(578).
p(580) :- p(579), q(580).
q(580) :- p(579), q(579).
p(581) :- p(580), q(581).
q(581) :- p(580), q(580).
p(582) :- p(581), q(582).
q(582) :- p(581), q(581).
p(583) :- p(582), q(583).
q(583) :- p(582), q(582).
p(584) :- p(583), q(584).
q(584) :- p(583), q(583).
p(585) :- p(584), q(585).
q(585) :- p(584), q(584).
p(586) :- p(585), q(586).
q(586) :- p(585), q(585).
p(587) :- p(586), q(587).
q(587) :- p(586), q(586).
p(588) :- p(587), q(588).
q(588) :- p(587), q(587).
p(589) :- p(588), q(589).
q(589) :- p(588), q(588).
p(590) :- p(589), q(590).
q(590) :- p(589), q(589).
p(591) :- p(590), q(591).
q(591) :- p(590), q(590).
p(592) :- p(591), q(592).
q(592) :- p(591), q(591).
p(593) :- p(592), q(593).
q(593) :- p(592), q(592).
p(594) :- p(593), q(594).
q(594) :- p(593), q(593).
p(595) :- p(594), q(595).
q(595) :- p(594), q(594).
p(596) :- p(595), q(596).
q(596) :- p(595), q(595).
p(597) :- p(596), q(597).
q(597) :- p(596), q(596).
p(598) :- p(597), q(598).
q(598) :- p(597), q(597).
p(599) :- p(598), q(599).
q(599) :- p(598), q(598).
p(600) :- p(599), q(600).
q(600) :- p(599), q(599).
p(601) :- p(600), q(601).
q(601) :- p(600), q(600).
p(602) :- p(601), q(602).
q(602) :- p(601), q(601).
p(603) :- p(602), q(603).
q(603) :- p(602), q(602).
p(604) :- p(603), q(604).
q(604) :- p(603), q(603).
p(605) :- p(604), q(605).
q(605) :- p(604), q(604).
p(606) :- p(605), q(606).
q(606) :- p(605), q(605).
p(607) :- p(606), q(607).
q(607) :- p(606), q(606).
p(608) :- p(607), q(608).
q(608) :- p(607), q(607).
p(609) :- p(608), q(609).
q(609) :- p(608), q(608).
p(610) :- p(609), q(610).
q(610) :- p(609), q(609).
p(611) :- p(610), q(611).
q(611) :- p(610), q(610).
p(612) :- p(611), q(612).
q(612) :- p(611), q(611).
p(613) :- p(612), q(613).
q(613) :- p(612), q(612).
p(614) :- p(613), q(614).
q(614) :- p(613), q(613).
p(615) :- p(614), q(615).
q(615) :- p(614), q(614).
p(616) :- p(615), q(616).
q(616) :- p(615), q(615).
p(617) :- p(616), q(617).
q(617) :- p(616), q(616).
p(618) :- p(617), q(618).
q(618) :- p(617), q(617).
p(619) :- p(618), q(619).
q(619) :- p(618), q(618).
p(620) :- p(619), q(620).
q(620) :- p(619), q(619).
p(621) :- p(620), q(621).
q(621) :- p(620), q(620).
p(622) :- p(621), q(622).
q(622) :- p(621), q(621).
p(623) :- p(622), q(623).
q(623) :- p(622), q(622).
p(624) :- p(623), q(624).
q(624) :- p(623), q(623).
p(625) :- p(624), q(625).
q(625) :- p(624), q(624).
p(626) :- p(625), q(626).
q(626) :- p(625), q(625).
p(627) :- p(626), q(627).
q(627) :- p(626), q(626).
p(628) :- p(627), q(628).
q(628) :- p(627), q(627).
p(629) :- p(628), q(629).
q(629) :- p(628), q(628).
p(630) :- p(629), q(630).
q(630) :- p(629), q(629).
p(631) :- p(630), q(631).
q(631) :- p(630), q(630).
p(632) :- p(631), q(632).
q(632) :- p(631), q(631).
p(633) :- p(632), q(633).
q(633) :- p(632), q(632).
p(634) :- p(633), q(634).
q(634) :- p(633), q(633).
p(635) :- p(634), q(635).
q(635) :- p(634), q(634).
p(636) :- p(635), q(636).
q(636) :- p(635), q(635).
p(637) :- p(636), q(637).
q(637) :- p(636), q(636).
p(638) :- p(637), q(638).
q(638) :- p(637), q(637).
p(639) :- p(638), q(639).
q(639) :- p(638), q(638).
p(640) :- p(639), q(640).
q(640) :- p(639), q(639).
p(641) :- p(640), q(641).
q(641) :- p(640), q(640).
p(642) :- p(641), q(642).
q(642) :- p(641), q(641).
p(643) :- p(642), q(643).
q(643) :- p(642), q(642).
p(644) :- p(643), q(644).
q(644) :- p(643), q(643).
p(645) :- p(644), q(645).
q(645) :- p(644), q(644).
p(646) :- p(645), q(646).
q(646) :- p(645), q(645).
p(647) :- p(646), q(647).
q(647) :- p(646), q(646).
p(648) :- p(647), q(648).
q(648) :- p(647), q(647).
p(649) :- p(648), q(649).
q(649) :- p(648), q(648).
p(650) :- p(649), q(650).
q(650) :- p(649), q(649).
p(651) :- p(650), q(651).
q(651) :- p(650), q(650).
p(652) :- p(651), q(652).
q(652) :- p(651), q(651).
p(653) :- p(652), q(653).
q(653) :- p(652), q(652).
p(654) :- p(653), q(654).
q(654) :- p(653), q(653).
p(655) :- p(654), q(655).
q(655) :- p(654), q(654).
p(656) :- p(655), q(656).
q(656) :- p(655), q(655).
p(657) :- p(656), q(657).
q(657) :- p(656), q(656).
p(658) :- p(657), q(658).
q(658) :- p(657), q(657).
p(659) :- p(658), q(659).
q(659) :- p(658), q(658).
p(660) :- p(659), q(660).
q(660) :- p(659), q(659).
p(661) :- p(660), q(661).
q(661) :- p(660), q(660).
p(662) :- p(661), q(662).
q(662) :- p(661), q(661).
p(663) :- p(662), q(663).
q(663) :- p(662), q(662).
p(664) :- p(663), q(664).
q(664) :- p(663), q(663).
p(665) :- p(664), q(665).
q(665) :- p(664), q(664).
p(666) :- p(665), q(666).
q(666) :- p(665), q(665).
p(667) :- p(666), q(667).
q(667) :- p(666), q(666).
p(668) :- p(667), q(668).
q(668) :- p(667), q(667).
p(669) :- p(668), q(669).
q(669) :- p(668), q(668).
p(670) :- p(669), q(670).
q(670) :- p(669), q(669).
p(671) :- p(670), q(671).
q(671) :- p(670), q(670).
p(672) :- p(671), q(672).
q(672) :- p(671), q(671).
p(673) :- p(672), q(673).
q(673) :- p(672), q(672).
p(674) :- p(673), q(674).
q(674) :- p(673), q(673).
p(675) :- p(674), q(675).
q(675) :- p(674), q(674).
p(676) :- p(675), q(676).
q(676) :- p(675), q(675).
p(677) :- p(676), q(677).
q(677) :- p(676), q(676).
p(678) :- p(677), q(678).
q(678) :- p(677), q(677).
p(679) :- p(678), q(679).
q(679) :- p(678), q(678).
p(680) :- p(679), q(680).
q(680) :- p(679), q(679).
p(681) :- p(680), q(681).
q(681) :- p(680), q(680).
p(682) :- p(681), q(682).
q(682) :- p(681), q(681).
p(683) :- p(682), q(683).
q(683) :- p(682), q(682).
p(684) :- p(683), q(684).
q(684) :- p(683), q(683).
p(685) :- p(684), q(685).
q(685) :- p(684), q(684).
p(686) :- p(685), q(686).
q(686) :- p(685), q(685).
p(687) :- p(686), q(687).
q(687) :- p(686), q(686).
p(688) :- p(687), q(688).
q(688) :- p(687), q(687).
p(689) :- p(688), q(689).
q(689) :- p(688), q(688).
p(690) :- p(689), q(690).
q(690) :- p(689), q(689).
p(691) :- p(690), q(691).
q(691) :- p(690), q(690).
p(692) :- p(691), q(692).
q(692) :- p(691), q(691).
p(693) :- p(692), q(693).
q(693) :- p(692), q(692).
p(694) :- p(693), q(694).
q(694) :- p(693), q(693).
p(695) :- p(694), q(695).
q(695) :- p(694), q(694).
p(696) :- p(695), q(696).
q(696) :- p(695), q(695).
p(697) :- p(696), q(697).
q(697) :- p(696), q(696).
p(698) :- p(697), q(698).
q(698) :- p(697), q(697).
p(699) :- p(698), q(699).
q(699) :- p(698), q(698).
p(700) :- p(699), q(700).
q(700) :- p(699), q(699).
p(701) :- p(700), q(701).
q(701) :- p(700), q(700).
p(702) :- p(701), q(702).
q(702) :- p(701), q(701).
p(703) :- p(702), q(703).
q(703) :- p(702), q(702).
p(704) :- p(703), q(704).
q(704) :- p(703), q(703).
p(705) :- p(704), q(705).
q(705) :- p(704), q(704).
p(706) :- p(705), q(706).
q(706) :- p(705), q(705).
p(707) :- p(706), q(707).
q(707) :- p(706), q(706).
p(708) :- p(707), q(708).
q(708) :- p(707), q(707).
p(709) :- p(708), q(709).
q(709) :- p(708), q(708).
p(710) :- p(709), q(710).
q(710) :- p(709), q(709).
p(711) :- p(710), q(711).
q(711) :- p(710), q(710).
p(712) :- p(711), q(712).
q(712) :- p(711), q(711).
p(713) :- p(712), q(713).
q(713) :- p(712), q(712).
p(714) :- p(713), q(714).
q(714) :- p(713), q(713).
p(715) :- p(714), q(715).
q(715) :- p(714), q(714).
p(716) :- p(715), q(716).
q(716) :- p(715), q(715).
p(717) :- p(716), q(717).
q(717) :- p(716), q(716).
p(718) :- p(717), q(718).
q(718) :- p(717), q(717).
p(719) :- p(718), q(719).
q(719) :- p(718), q(718).
p(720) :- p(719), q(720).
q(720) :- p(719), q(719).
p(721) :- p(720), q(721).
q(721) :- p(720), q(720).
p(722) :- p(721), q(722).
q(722) :- p(721), q(721).
p(723) :- p(722), q(723).
q(723) :- p(722), q(722).
p(724) :- p(723), q(724).
q(724) :- p(723), q(723).
p(725) :- p(724), q(725).
q(725) :- p(724), q(724).
p(726) :- p(725), q(726).
q(726) :- p(725), q(725).
p(727) :- p(726), q(727).
q(727) :- p(726), q(726).
p(728) :- p(727), q(728).
q(728) :- p(727), q(727).
p(729) :- p(728), q(729).
q(729) :- p(728), q(728).
p(730) :- p(729), q(730).
q(730) :- p(729), q(729).
p(731) :- p(730), q(731).
q(731) :- p(730), q(730).
p(732) :- p(731), q(732).
q(732) :- p(731), q(731).
p(733) :- p(732), q(733).
q(733) :- p(732), q(732).
p(734) :- p(733), q(734).
q(734) :- p(733), q(733).
p(735) :- p(734), q(735).
q(735) :- p(734), q(734).
p(736) :- p(735), q(736).
q(736) :- p(735), q(735).
p(737) :- p(736), q(737).
q(737) :- p(736), q(736).
p(738) :- p(737), q(738).
q(738) :- p(737), q(737).
p(739) :- p(738), q(739).
q(739) :- p(738), q(738).
p(740) :- p(739), q(740).
q(740) :- p(739), q(739).
p(741) :- p(740), q(741).
q(741) :- p(740), q(740).
p(742) :- p(741), q(742).
q(742) :- p(741), q(741).
p(743) :- p(742), q(743).
q(743) :- p(742), q(742).
p(744) :- p(743), q(744).
q(744) :- p(743), q(743).
p(745) :- p(744), q(745).
q(745) :- p(744), q(744).
p(746) :- p(745), q(746).
q(746) :- p(745), q(745).
p(747) :- p(746), q(747).
q(747) :- p(746), q(746).
p(748) :- p(747), q(748).
q(748) :- p(747), q(747).
p(749) :- p(748), q(749).
q(749) :- p(748), q(748).
p(750) :- p(749), q(750).
q(750) :- p(749), q(749).
p(751) :- p(750), q(751).
q(751) :- p(750), q(750).
p(752) :- p(751), q(752).
q(752) :- p(751), q(751).
p(753) :- p(752), q(753).
q(753) :- p(752), q(752).
p(754) :- p(753), q(754).
q(754) :- p(753), q(753).
p(755) :- p(754), q(755).
q(755) :- p(754), q(754).
p(756) :- p(755), q(756).
q(756) :- p(755), q(755).
p(757) :- p(756), q(757).
q(757) :- p(756), q(756).
p(758) :- p(757), q(758).
q(758) :- p(757), q(757).
p(759) :- p(758), q(759).
q(759) :- p(758), q(758).
p(760) :- p(759), q(760).
q(760) :- p(759), q(759).
p(761) :- p(760), q(761).
q(761) :- p(760), q(760).
p(762) :- p(761), q(762).
q(762) :- p(761), q(761).
p(763) :- p(762), q(763).
q(763) :- p(762), q(762).
p(764) :- p(763), q(764).
q(764) :- p(763), q(763).
p(765) :- p(764), q(765).
q(765) :- p(764), q(764).
p(766) :- p(765), q(766).
q(766) :- p(765), q(765).
p(767) :- p(766), q(767).
q(767) :- p(766), q(766).
p(768) :- p(767), q(768).
q(768) :- p(767), q(767).
p(769) :- p(768), q(769).
q(769) :- p(768), q(768).
p(770) :- p(769), q(770).
q(770) :- p(769), q(769).
p(771) :- p(770), q(771).
q(771) :- p(770), q(770).
p(772) :- p(771), q(772).
q(772) :- p(771), q(771).
p(773) :- p(772), q(773).
q(773) :- p(772), q(772).
p(774) :- p(773), q(774).
q(774) :- p(773), q(773).
p(775) :- p(774), q(775).
q(775) :- p(774), q(774).
p(776) :- p(775), q(776).
q(776) :- p(775), q(775).
p(777) :- p(776), q(777).
q(777) :- p(776), q(776).
p(778) :- p(777), q(778).
q(778) :- p(777), q(777).
p(779) :- p(778), q(779).
q(779) :- p(778), q(778).
p(780) :- p(779), q(780).
q(780) :- p(779), q(779).
p(781) :- p(780), q(781).
q(781) :- p(780), q(780).
p(782) :- p(781), q(782).
q(782) :- p(781), q(781).
p(783) :- p(782), q(783).
q(783) :- p(782), q(782).
p(784) :- p(783), q(784).
q(784) :- p(783), q(783).
p(785) :- p(784), q(785).
q(785) :- p(784), q(784).
p(786) :- p(785), q(786).
q(786) :- p(785), q(785).
p(787) :- p(786), q(787).
q(787) :- p(786), q(786).
p(788) :- p(787), q(788).
q(788) :- p(787), q(787).
p(789) :- p(788), q(789).
q(789) :- p(788), q(788).
p(790) :- p(789), q(790).
q(790) :- p(789), q(789).
p(791) :- p(790), q(791).
q(791) :- p(790), q(790).
p(792) :- p(791), q(792).
q(792) :- p(791), q(791).
p(793) :- p(792), q(793).
q(793) :- p(792), q(792).
p(794) :- p(793), q(794).
q(794) :- p(793), q(793).
p(795) :- p(794), q(795).
q(795) :- p(794), q(794).
p(796) :- p(795), q(796).
q(796) :- p(795), q(795).
p(797) :- p(796), q(797).
q(797) :- p(796), q(796).
p(798) :- p(797), q(798).
q(798) :- p(797), q(797).
p(799) :- p(798), q(799).
q(799) :- p(798), q(798).
p(800) :- p(799), q(800).
q(800) :- p(799), q(799).
p(801) :- p(800), q(801).
q(801) :- p(800), q(800).
p(802) :- p(801), q(802).
q(802) :- p(801), q(801).
p(803) :- p(802), q(803).
q(803) :- p(802), q(802).
p(804) :- p(803), q(804).
q(804) :- p(803), q(803).
p(805) :- p(804), q(805).
q(805) :- p(804), q(804).
p(806) :- p(805), q(806).
q(806) :- p(805), q(805).
p(807) :- p(806), q(807).
q(807) :- p(806), q(806).
p(808) :- p(807), q(808).
q(808) :- p(807), q(807).
p(809) :- p(808), q(809).
q(809) :- p(808), q(808).
p(810) :- p(809), q(810).
q(810) :- p(809), q(809).
p(811) :- p(810), q(811).
q(811) :- p(810), q(810).
p(812) :- p(811), q(812).
q(812) :- p(811), q(811).
p(813) :- p(812), q(813).
q(813) :- p(812), q(812).
p(814) :- p(813), q(814).
q(814) :- p(813), q(813).
p(815) :- p(814), q(815).
q(815) :- p(814), q(814).
p(816) :- p(815), q(816).
q(816) :- p(815), q(815).
p(817) :- p(816), q(817).
q(817) :- p(816), q(816).
p(818) :- p(817), q(818).
q(818) :- p(817), q(817).
p(819) :- p(818), q(819).
q(819) :- p(818), q(818).
p(820) :- p(819), q(820).
q(820) :- p(819), q(819).
p(821) :- p(820), q(821).
q(821) :- p(820), q(820).
p(822) :- p(821), q(822).
q(822) :- p(821), q(821).
p(823) :- p(822), q(823).
q(823) :- p(822), q(822).
p(824) :- p(823), q(824).
q(824) :- p(823), q(823).
p(825) :- p(824), q(825).
q(825) :- p(824), q(824).
p(826) :- p(825), q(826).
q(826) :- p(825), q(825).
p(827) :- p(826), q(827).
q(827) :- p(826), q(826).
p(828) :- p(827), q(828).
q(828) :- p(827), q(827).
p(829) :- p(828), q(829).
q(829) :- p(828), q(828).
p(830) :- p(829), q(830).
q(830) :- p(829), q(829).
p(831) :- p(830), q(831).
q(831) :- p(830), q(830).
p(832) :- p(831), q(832).
q(832) :- p(831), q(831).
p(833) :- p(832), q(833).
q(833) :- p(832), q(832).
p(834) :- p(833), q(834).
q(834) :- p(833), q(833).
p(835) :- p(834), q(835).
q(835) :- p(834), q(834).
p(836) :- p(835), q(836).
q(836) :- p(835), q(835).
p(837) :- p(836), q(837).
q(837) :- p(836), q(836).
p(838) :- p(837), q(838).
q(838) :- p(837), q(837).
p(839) :- p(838), q(839).
q(839) :- p(838), q(838).
p(840) :- p(839), q(840).
q(840) :- p(839), q(839).
p(841) :- p(840), q(841).
q(841) :- p(840), q(840).
p(842) :- p(841), q(842).
q(842) :- p(841), q(841).
p(843) :- p(842), q(843).
q(843) :- p(842), q(842).
p(844) :- p(843), q(844).
q(844) :- p(843), q(843).
p(845) :- p(844), q(845).
q(845) :- p(844), q(844).
p(846) :- p(845), q(846).
q(846) :- p(845), q(845).
p(847) :- p(846), q(847).
q(847) :- p(846), q(846).
p(848) :- p(847), q(848).
q(848) :- p(847), q(847).
p(849) :- p(848), q(849).
q(849) :- p(848), q(848).
p(850) :- p(849), q(850).
q(850) :- p(849), q(849).
p(851) :- p(850), q(851).
q(851) :- p(850), q(850).
p(852) :- p(851), q(852).
q(852) :- p(851), q(851).
p(853) :- p(852), q(853).
q(853) :- p(852), q(852).
p(854) :- p(853), q(854).
q(854) :- p(853), q(853).
p(855) :- p(854), q(855).
q(855) :- p(854), q(854).
p(856) :- p(855), q(856).
q(856) :- p(855), q(855).
p(857) :- p(856), q(857).
q(857) :- p(856), q(856).
p(858) :- p(857), q(858).
q(858) :- p(857), q(857).
p(859) :- p(858), q(859).
q(859) :- p(858), q(858).
p(860) :- p(859), q(860).
q(860) :- p(859), q(859).
p(861) :- p(860), q(861).
q(861) :- p(860), q(860).
p(862) :- p(861), q(862).
q(862) :- p(861), q(861).
p(863) :- p(862), q(863).
q(863) :- p(862), q(862).
p(864) :- p(863), q(864).
q(864) :- p(863), q(863).
p(865) :- p(864), q(865).
q(865) :- p(864), q(864).
p(866) :- p(865), q(866).
q(866) :- p(865), q(865).
p(867) :- p(866), q(867).
q(867) :- p(866), q(866).
p(868) :- p(867), q(868).
q(868) :- p(867), q(867).
p(869) :- p(868), q(869).
q(869) :- p(868), q(868).
p(870) :- p(869), q(870).
q(870) :- p(869), q(869).
p(871) :- p(870), q(871).
q(871) :- p(870), q(870).
p(872) :- p(871), q(872).
q(872) :- p(871), q(871).
p(873) :- p(872), q(873).
q(873) :- p(872), q(872).
p(874) :- p(873), q(874).
q(874) :- p(873), q(873).
p(875) :- p(874), q(875).
q(875) :- p(874), q(874).
p(876) :- p(875), q(876).
q(876) :- p(875), q(875).
p(877) :- p(876), q(877).
q(877) :- p(876), q(876).
p(878) :- p(877), q(878).
q(878) :- p(877), q(877).
p(879) :- p(878), q(879).
q(879) :- p(878), q(878).
p(880) :- p(879), q(880).
q(880) :- p(879), q(879).
p(881) :- p(880), q(881).
q(881) :- p(880), q(880).
p(882) :- p(881), q(882).
q(882) :- p(881), q(881).
p(883) :- p(882), q(883).
q(883) :- p(882), q(882).
p(884) :- p(883), q(884).
q(884) :- p(883), q(883).
p(885) :- p(884), q(885).
q(885) :- p(884), q(884).
p(886) :- p(885), q(886).
q(886) :- p(885), q(885).
p(887) :- p(886), q(887).
q(887) :- p(886), q(886).
p(888) :- p(887), q(888).
q(888) :- p(887), q(887).
p(889) :- p(888), q(889).
q(889) :- p(888), q(888).
p(890) :- p(889), q(890).
q(890) :- p(889), q(889).
p(891) :- p(890), q(891).
q(891) :- p(890), q(890).
p(892) :- p(891), q(892).
q(892) :- p(891), q(891).
p(893) :- p(892), q(893).
q(893) :- p(892), q(892).
p(894) :- p(893), q(894).
q(894) :- p(893), q(893).
p(895) :- p(894), q(895).
q(895) :- p(894), q(894).
p(896) :- p(895), q(896).
q(896) :- p(895), q(895).
p(897) :- p(896), q(897).
q(897) :- p(896), q(896).
p(898) :- p(897), q(898).
q(898) :- p(897), q(897).
p(899) :- p(898), q(899).
q(899) :- p(898), q(898).
p(900) :- p(899), q(900).
q(900) :- p(899), q(899).
p(901) :- p(900), q(901).
q(901) :- p(900), q(900).
p(902) :- p(901), q(902).
q(902) :- p(901), q(901).
p(903) :- p(902), q(903).
q(903) :- p(902), q(902).
p(904) :- p(903), q(904).
q(904) :- p(903), q(903).
p(905) :- p(904), q(905).
q(905) :- p(904), q(904).
p(906) :- p(905), q(906).
q(906) :- p(905), q(905).
p(907) :- p(906), q(907).
q(907) :- p(906), q(906).
p(908) :- p(907), q(908).
q(908) :- p(907), q(907).
p(909) :- p(908), q(909).
q(909) :- p(908), q(908).
p(910) :- p(909), q(910).
q(910) :- p(909), q(909).
p(911) :- p(910), q(911).
q(911) :- p(910), q(910).
p(912) :- p(911), q(912).
q(912) :- p(911), q(911).
p(913) :- p(912), q(913).
q(913) :- p(912), q(912).
p(914) :- p(913), q(914).
q(914) :- p(913), q(913).
p(915) :- p(914), q(915).
q(915) :- p(914), q(914).
p(916) :- p(915), q(916).
q(916) :- p(915), q(915).
p(917) :- p(916), q(917).
q(917) :- p(916), q(916).
p(918) :- p(917), q(918).
q(918) :- p(917), q(917).
p(919) :- p(918), q(919).
q(919) :- p(918), q(918).
p(920) :- p(919), q(920).
q(920) :- p(919), q(919).
p(921) :- p(920), q(921).
q(921) :- p(920), q(920).
p(922) :- p(921), q(922).
q(922) :- p(921), q(921).
p(923) :- p(922), q(923).
q(923) :- p(922), q(922).
p(924) :- p(923), q(924).
q(924) :- p(923), q(923).
p(925) :- p(924), q(925).
q(925) :- p(924), q(924).
p(926) :- p(925), q(926).
q(926) :- p(925), q(925).
p(927) :- p(926), q(927).
q(927) :- p(926), q(926).
p(928) :- p(927), q(928).
q(928) :- p(927), q(927).
p(929) :- p(928), q(929).
q(929) :- p(928), q(928).
p(930) :- p(929), q(930).
q(930) :- p(929), q(929).
p(931) :- p(930), q(931).
q(931) :- p(930), q(930).
p(932) :- p(931), q(932).
q(932) :- p(931), q(931).
p(933) :- p(932), q(933).
q(933) :- p(932), q(932).
p(934) :- p(933), q(934).
q(934) :- p(933), q(933).
p(935) :- p(934), q(935).
q(935) :- p(934), q(934).
p(936) :- p(935), q(936).
q(936) :- p(935), q(935).
p(937) :- p(936), q(937).
q(937) :- p(936), q(936).
p(938) :- p(937), q(938).
q(938) :- p(937), q(937).
p(939) :- p(938), q(939).
q(939) :- p(938), q(938).
p(940) :- p(939), q(940).
q(940) :- p(939), q(939).
p(941) :- p(940), q(941).
q(941) :- p(940), q(940).
p(942) :- p(941), q(942).
q(942) :- p(941), q(941).
p(943) :- p(942), q(943).
q(943) :- p(942), q(942).
p(944) :- p(943), q(944).
q(944) :- p(943), q(943).
p(945) :- p(944), q(945).
q(945) :- p(944), q(944).
p(946) :- p(945), q(946).
q(946) :- p(945), q(945).
p(947) :- p(946), q(947).
q(947) :- p(946), q(946).
p(948) :- p(947), q(948).
q(948) :- p(947), q(947).
p(949) :- p(948), q(949).
q(949) :- p(948), q(948).
p(950) :- p(949), q(950).
q(950) :- p(949), q(949).
p(951) :- p(950), q(951).
q(951) :- p(950), q(950).
p(952) :- p(951), q(952).
q(952) :- p(951), q(951).
p(953) :- p(952), q(953).
q(953) :- p(952), q(952).
p(954) :- p(953), q(954).
q(954) :- p(953), q(953).
p(955) :- p(954), q(955).
q(955) :- p(954), q(954).
p(956) :- p(955), q(956).
q(956) :- p(955), q(955).
p(957) :- p(956), q(957).
q(957) :- p(956), q(956).
p(958) :- p(957), q(958).
q(958) :- p(957), q(957).
p(959) :- p(958), q(959).
q(959) :- p(958), q(958).
p(960) :- p(959), q(960).
q(960) :- p(959), q(959).
p(961) :- p(960), q(961).
q(961) :- p(960), q(960).
p(962) :- p(961), q(962).
q(962) :- p(961), q(961).
p(963) :- p(962), q(963).
q(963) :- p(962), q(962).
p(964) :- p(963), q(964).
q(964) :- p(963), q(963).
p(965) :- p(964), q(965).
q(965) :- p(964), q(964).
p(966) :- p(965), q(966).
q(966) :- p(965), q(965).
p(967) :- p(966), q(967).
q(967) :- p(966), q(966).
p(968) :- p(967), q(968).
q(968) :- p(967), q(967).
p(969) :- p(968), q(969).
q(969) :- p(968), q(968).
p(970) :- p(969), q(970).
q(970) :- p(969), q(969).
p(971) :- p(970), q(971).
q(971) :- p(970), q(970).
p(972) :- p(971), q(972).
q(972) :- p(971), q(971).
p(973) :- p(972), q(973).
q(973) :- p(972), q(972).
p(974) :- p(973), q(974).
q(974) :- p(973), q(973).
p(975) :- p(974), q(975).
q(975) :- p(974), q(974).
p(976) :- p(975), q(976).
q(976) :- p(975), q(975).
p(977) :- p(976), q(977).
q(977) :- p(976), q(976).
p(978) :- p(977), q(978).
q(978) :- p(977), q(977).
p(979) :- p(978), q(979).
q(979) :- p(978), q(978).
p(980) :- p(979), q(980).
q(980) :- p(979), q(979).
p(981) :- p(980), q(981).
q(981) :- p(980), q(980).
p(982) :- p(981), q(982).
q(982) :- p(981), q(981).
p(983) :- p(982), q(983).
q(983) :- p(982), q(982).
p(984) :- p(983), q(984).
q(984) :- p(983), q(983).
p(985) :- p(984), q(985).
q(985) :- p(984), q(984).
p(986) :- p(985), q(986).
q(986) :- p(985), q(985).
p(987) :- p(986), q(987).
q(987) :- p(986), q(986).
p(988) :- p(987), q(988).
q(988) :- p(987), q(987).
p(989) :- p(988), q(989).
q(989) :- p(988), q(988).
p(990) :- p(989), q(990).
q(990) :- p(989), q(989).
p(991) :- p(990), q(991).
q(991) :- p(990), q(990).
p(992) :- p(991), q(992).
q(992) :- p(991), q(991).
p(993) :- p(992), q(993).
q(993) :- p(992), q(992).
p(994) :- p(993), q(994).
q(994) :- p(993), q(993).
p(995) :- p(994), q(995).
q(995) :- p(994), q(994).
p(996) :- p(995), q(996).
q(996) :- p(995), q(995).
p(997) :- p(996), q(997).
q(997) :- p(996), q(996).
p(998) :- p(997), q(998).
q(998) :- p(997), q(997).
p(999) :- p(998), q(999).
q(999) :- p(998), q(998).
p(1000) :- p(999), q(1000).
q(1000) :- p(999), q(999).