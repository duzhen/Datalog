p(0).

p(1) :- not p(0).
p(1) :- p(0).