person(ann).
person(bertrand).
person(charles).
person(dorothy).
person(evelyn).
person(fred).
person(george).
person(hilary).
par(dorothy, george).
par(evelyn, george).
par(bertrand, dorothy).
par(ann, dorothy).
par(ann, hilary).
par(charles, evelyn).

sgc(X, X) :- person(X).
sgc(X, Y) :- par(X, X1), sgc(X1, Y1), par(Y, Y1).

sgc(ann, dorothy)?
sgc(ann, charles)?
