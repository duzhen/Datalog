e(a,b,1).
e(b,c,1).
e(a,c,1).
e(c,d,1).
e(d,e,1).
e(c,e,1).
e(a,f,1).
e(f,e,1).

c(1, 1, 1).
c(2, 1, 2).
c(3, 1, 3).
c(4, 1, 4).
c(2, 2, 1).
c(4, 2, 2).
c(6, 2, 3).
c(8, 2, 4).
c(3, 3, 1).
c(6, 3, 2).
c(9, 3, 3).
c(12, 3, 4).
c(4, 4, 1).
c(8, 4, 2).
c(12, 4, 3).
c(16, 4, 4).

c1(2, 1, 1).
c1(3, 1, 2).
c1(4, 1, 3).
c1(5, 1, 4).
c1(3, 2, 1).
c1(5, 2, 2).
c1(7, 2, 3).
c1(9, 2, 4).
c1(4, 3, 1).
c1(7, 3, 2).
c1(10, 3, 3).
c1(13, 3, 4).
c1(5, 4, 1).
c1(9, 4, 2).
c1(13, 4, 3).
c1(17, 4, 4).

p(X, Y, N) :- e(X, Y, N).
p(X, Y, N) :- p(X, Z, N1), p(Z, Y, N2), c(N, N1, N2).
p(X, Y, N) :- p(X, Y, N0), p(X, Z, N1), p(Z, Y, N2), c1(N, N1, N2).

p(a, e, N)?
