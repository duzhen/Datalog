parent(alice, bob).
parent(alice, bill).
parent(bob, carol).
parent(carol, dennis).
parent(carol, david).
age(alice, 30.00).
age(bob, 40.500).
weight(bob, 10056.7000).

ancestor(X, Y) :- parent(X, Y).
ancestor(X, Y) :- ancestor(X, Z), ancestor(Z, Y).
family(X, Y) :- ancestor(X, Y).
family(X, Y) :- family(Y, X).

details(X, Age, Address, Weight) :- age(X, Age), address(X, Address), weight(X, Weight).
details(bob, Age, Address, Weight)?


age(alice, Age)?
age(bob, Age)?
weight(bob, Weight)?
family(X, Y)?
family(alice, Y)?
family(alex, Y)?
ancestor(bob, Y)?

address(bob, Address)?
address(carol, Address)?