p(0).

k(1) :- not q(0).
q(0) :- not p(1).
% p->q->k

q(X)?
k(X)?