edge(a, b).
edge(a, c).
edge(b, d).
edge(c, d).
edge(1, 2).
not edge(f, e).

path(X, Y) :- edge(X, Y), X==Y.
path(X, Y) :- path(X, Z), path(Z, Y).
path(X, X) :- not edge(X, X).

path(a, b)?
path(f, X), V == e?
path(a, X), path(X, d)?
not path(f, e)?